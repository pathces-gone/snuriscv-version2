module snurisc(
    input i_reset,
    input i_clk,
    input i_clock_en
    );

    // TODO
endmodule