/*
* Module : snurisc_core
* Author : Evan.Park
* Date   : May 29, 2023
* Description: This module is snurisc-core module, which is fabricated Datapath and control-logic.
*/
`timescale 1ns / 1ps