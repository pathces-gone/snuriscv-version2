/*
* Module : snurisc_top
* Author : Evan.Park
* Date   : May 29, 2023
* Description: This module is snurisc-top module, which is System-on-chip
*              fabricating I$, D$, snurisc-core, ... 
*/
`timescale 1ns / 1ps

module snurisc(
    input i_reset,
    input i_clk,
    input i_clock_en
    );

    // TODO
endmodule